
`define UIO_OE_INPUT   1'b0
`define UIO_OE_OUTPUT  1'b1
